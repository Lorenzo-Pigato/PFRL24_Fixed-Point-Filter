library ieee;
use ieee.std_logic_1164.all;

entity CLOCK_GATE is
end clockgate;

architecture clockgate of clockgate is
	port(
			EN			:	in std_logic;
			CLK		:	in std_logic;
			CLK		:	out std_logic;
			NOT_CLK	:	out std_logic
		);
begin


end CLOCK_GATE;

